module Adder(
    input [2:0] A,
    input [2:0] B,
    output [2:0] result
    );
    assign result = A + B;
endmodule
